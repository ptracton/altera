// testing_tb.v

// Generated using ACDS version 13.1 162 at 2014.06.02.17:44:15

`timescale 1 ps / 1 ps
module testing_tb (
	);

	wire        testing_inst_clk_bfm_clk_clk;                   // testing_inst_clk_bfm:clk -> [testing_inst:clk_clk, testing_inst_reset_bfm:clk]
	wire        testing_inst_reset_bfm_reset_reset;             // testing_inst_reset_bfm:reset -> testing_inst:reset_reset_n
	wire  [7:0] testing_inst_leds_output_export;                // testing_inst:leds_output_export -> testing_inst_leds_output_bfm:sig_export
	wire  [7:0] testing_inst_switches_input_bfm_conduit_export; // testing_inst_switches_input_bfm:sig_export -> testing_inst:switches_input_export

	testing testing_inst (
		.clk_clk               (testing_inst_clk_bfm_clk_clk),                   //            clk.clk
		.reset_reset_n         (testing_inst_reset_bfm_reset_reset),             //          reset.reset_n
		.leds_output_export    (testing_inst_leds_output_export),                //    leds_output.export
		.switches_input_export (testing_inst_switches_input_bfm_conduit_export)  // switches_input.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) testing_inst_clk_bfm (
		.clk (testing_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) testing_inst_reset_bfm (
		.reset (testing_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (testing_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm testing_inst_leds_output_bfm (
		.sig_export (testing_inst_leds_output_export)  // conduit.export
	);

	altera_conduit_bfm_0002 testing_inst_switches_input_bfm (
		.sig_export (testing_inst_switches_input_bfm_conduit_export)  // conduit.export
	);

endmodule
