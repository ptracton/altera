module top();
   pattern_generator_tb tb();
   test_program pgm();
endmodule