// interrupt_example_tb.v

// Generated using ACDS version 13.1 162 at 2014.06.06.12:54:28

`timescale 1 ps / 1 ps
module interrupt_example_tb (
			     );

   wire        interrupt_example_inst_clk_bfm_clk_clk;                   // interrupt_example_inst_clk_bfm:clk -> [interrupt_example_inst:clk_clk, interrupt_example_inst_reset_bfm:clk]
   wire        interrupt_example_inst_reset_bfm_reset_reset;             // interrupt_example_inst_reset_bfm:reset -> interrupt_example_inst:reset_reset_n
   reg [7:0]   interrupt_example_inst_switches_input_bfm_conduit_export; // interrupt_example_inst_switches_input_bfm:sig_export -> interrupt_example_inst:switches_input_export
   wire [7:0]  interrupt_example_inst_leds_output_export;                // interrupt_example_inst:leds_output_export -> interrupt_example_inst_leds_output_bfm:sig_export

   interrupt_example interrupt_example_inst (
					     .clk_clk               (interrupt_example_inst_clk_bfm_clk_clk),                   //            clk.clk
					     .reset_reset_n         (interrupt_example_inst_reset_bfm_reset_reset),             //          reset.reset_n
					     .switches_input_export (interrupt_example_inst_switches_input_bfm_conduit_export), // switches_input.export
					     .leds_output_export    (interrupt_example_inst_leds_output_export)                 //    leds_output.export
					     );

   altera_avalon_clock_source #(
				.CLOCK_RATE (50000000),
				.CLOCK_UNIT (1)
				) interrupt_example_inst_clk_bfm (
								  .clk (interrupt_example_inst_clk_bfm_clk_clk)  // clk.clk
								  );

   altera_avalon_reset_source #(
				.ASSERT_HIGH_RESET    (0),
				.INITIAL_RESET_CYCLES (50)
				) interrupt_example_inst_reset_bfm (
								    .reset (interrupt_example_inst_reset_bfm_reset_reset), // reset.reset_n
								    .clk   (interrupt_example_inst_clk_bfm_clk_clk)        //   clk.clk
								    );

/* -----\/----- EXCLUDED -----\/-----
   altera_conduit_bfm interrupt_example_inst_switches_input_bfm (
								 .sig_export (interrupt_example_inst_switches_input_bfm_conduit_export)  // conduit.export
								 );
 -----/\----- EXCLUDED -----/\----- */

   altera_conduit_bfm_0002 interrupt_example_inst_leds_output_bfm (
								   .sig_export (interrupt_example_inst_leds_output_export)  // conduit.export
								   );

   always @(posedge interrupt_example_inst_clk_bfm_clk_clk)
     if (!interrupt_example_inst_reset_bfm_reset_reset) begin
	interrupt_example_inst_switches_input_bfm_conduit_export <= 8'h00;	
     end else if (interrupt_example_inst_leds_output_export[0]) begin
	interrupt_example_inst_switches_input_bfm_conduit_export <= 8'h01;
     end else begin
	interrupt_example_inst_switches_input_bfm_conduit_export <= 8'h00;	
     end

endmodule
